** Layout Netlist, pvs precompare
** 

.subckt sarafe_nsw CLKB ENL0<0> ENL0<1> ENL0<2> ENL1<0> ENL1<1> ENL1<2> ENL2<0> ENL2<1> ENL2<2> ENL3<0> ENL3<1> ENL3<2> ENL4<0> ENL4<1> ENL4<2> ENL5<0> ENL5<1> ENL5<2> ENL6<0> 
+ ENL6<1> ENL6<2> ENL7<0> ENL7<1> ENL7<2> ENR0<0> ENR0<1> ENR0<2> ENR1<0> ENR1<1> ENR1<2> ENR2<0> ENR2<1> ENR2<2> ENR3<0> ENR3<1> ENR3<2> ENR4<0> ENR4<1> ENR4<2> 
+ ENR5<0> ENR5<1> ENR5<2> ENR6<0> ENR6<1> ENR6<2> ENR7<0> ENR7<1> ENR7<2> INM INP OSM OSP OUTM OUTP VDD VOL<0> VOL<1> VOL<2> VOL<3> 
+ VOL<4> VOL<5> VOL<6> VOL<7> VOR<0> VOR<1> VOR<2> VOR<3> VOR<4> VOR<5> VOR<6> VOR<7> VREF<0> VREF<1> VREF<2> VSS 
MX84/X99/X9/X14/X3/M0 X84/X99/X9/6 X84/X99/X9/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X9/X14/X4/M0 VSS X84/X99/X9/6 X84/X99/X9/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X9/X15/X3/M0 X84/X99/X9/7 X84/X99/X9/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X9/X15/X4/M0 VSS X84/X99/X9/7 X84/X99/X9/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X24/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X24/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X25/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X25/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X26/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X26/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X27/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X27/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X28/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X28/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X29/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X29/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X30/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X30/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X31/X3/M0 VOL<7> ENL7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X10/X31/X4/M0 VREF<0> ENL7<0> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X24/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X24/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X25/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X25/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X26/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X26/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X27/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X27/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X28/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X28/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X29/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X29/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X30/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X30/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X31/X3/M0 VOL<7> ENL7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X11/X31/X4/M0 VREF<1> ENL7<1> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X24/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X24/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X25/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X25/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X26/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X26/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X27/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X27/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X28/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X28/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X29/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X29/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X30/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X30/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X31/X3/M0 VOL<7> ENL7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X99/X12/X31/X4/M0 VREF<2> ENL7<2> VOL<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X12/X14/X3/M0 X84/X116/X12/6 X84/X116/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X12/X14/X4/M0 VSS X84/X116/X12/6 X84/X116/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X12/X15/X3/M0 X84/X116/X12/7 X84/X116/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X12/X15/X4/M0 VSS X84/X116/X12/7 X84/X116/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X13/X16/X3/M0 VOL<0> ENL0<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X13/X16/X4/M0 VREF<0> ENL0<0> VOL<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X13/X17/X3/M0 VOL<0> ENL0<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X13/X17/X4/M0 VREF<0> ENL0<0> VOL<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X14/X16/X3/M0 VOL<0> ENL0<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X14/X16/X4/M0 VREF<1> ENL0<1> VOL<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X14/X17/X3/M0 VOL<0> ENL0<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X14/X17/X4/M0 VREF<1> ENL0<1> VOL<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X15/X16/X3/M0 VOL<0> ENL0<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X15/X16/X4/M0 VREF<2> ENL0<2> VOL<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X15/X17/X3/M0 VOL<0> ENL0<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X116/X15/X17/X4/M0 VREF<2> ENL0<2> VOL<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X12/X14/X3/M0 X84/X117/X12/6 X84/X117/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X12/X14/X4/M0 VSS X84/X117/X12/6 X84/X117/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X12/X15/X3/M0 X84/X117/X12/7 X84/X117/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X12/X15/X4/M0 VSS X84/X117/X12/7 X84/X117/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X13/X16/X3/M0 VOL<2> ENL2<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X13/X16/X4/M0 VREF<0> ENL2<0> VOL<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X13/X17/X3/M0 VOL<2> ENL2<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X13/X17/X4/M0 VREF<0> ENL2<0> VOL<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X14/X16/X3/M0 VOL<2> ENL2<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X14/X16/X4/M0 VREF<1> ENL2<1> VOL<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X14/X17/X3/M0 VOL<2> ENL2<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X14/X17/X4/M0 VREF<1> ENL2<1> VOL<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X15/X16/X3/M0 VOL<2> ENL2<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X15/X16/X4/M0 VREF<2> ENL2<2> VOL<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X15/X17/X3/M0 VOL<2> ENL2<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X117/X15/X17/X4/M0 VREF<2> ENL2<2> VOL<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X12/X14/X3/M0 X84/X118/X12/6 X84/X118/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X12/X14/X4/M0 VSS X84/X118/X12/6 X84/X118/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X12/X15/X3/M0 X84/X118/X12/7 X84/X118/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X12/X15/X4/M0 VSS X84/X118/X12/7 X84/X118/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X13/X16/X3/M0 VOL<4> ENL4<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X13/X16/X4/M0 VREF<0> ENL4<0> VOL<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X13/X17/X3/M0 VOL<4> ENL4<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X13/X17/X4/M0 VREF<0> ENL4<0> VOL<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X14/X16/X3/M0 VOL<4> ENL4<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X14/X16/X4/M0 VREF<1> ENL4<1> VOL<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X14/X17/X3/M0 VOL<4> ENL4<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X14/X17/X4/M0 VREF<1> ENL4<1> VOL<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X15/X16/X3/M0 VOL<4> ENL4<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X15/X16/X4/M0 VREF<2> ENL4<2> VOL<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X15/X17/X3/M0 VOL<4> ENL4<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X118/X15/X17/X4/M0 VREF<2> ENL4<2> VOL<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X12/X14/X3/M0 X84/X119/X12/6 X84/X119/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X12/X14/X4/M0 VSS X84/X119/X12/6 X84/X119/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X12/X15/X3/M0 X84/X119/X12/7 X84/X119/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X12/X15/X4/M0 VSS X84/X119/X12/7 X84/X119/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X13/X16/X3/M0 VOL<1> ENL1<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X13/X16/X4/M0 VREF<0> ENL1<0> VOL<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X13/X17/X3/M0 VOL<1> ENL1<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X13/X17/X4/M0 VREF<0> ENL1<0> VOL<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X14/X16/X3/M0 VOL<1> ENL1<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X14/X16/X4/M0 VREF<1> ENL1<1> VOL<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X14/X17/X3/M0 VOL<1> ENL1<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X14/X17/X4/M0 VREF<1> ENL1<1> VOL<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X15/X16/X3/M0 VOL<1> ENL1<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X15/X16/X4/M0 VREF<2> ENL1<2> VOL<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X15/X17/X3/M0 VOL<1> ENL1<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X119/X15/X17/X4/M0 VREF<2> ENL1<2> VOL<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X12/X14/X3/M0 X84/X120/X12/6 X84/X120/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X12/X14/X4/M0 VSS X84/X120/X12/6 X84/X120/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X12/X15/X3/M0 X84/X120/X12/7 X84/X120/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X12/X15/X4/M0 VSS X84/X120/X12/7 X84/X120/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X13/X16/X3/M0 VOL<3> ENL3<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X13/X16/X4/M0 VREF<0> ENL3<0> VOL<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X13/X17/X3/M0 VOL<3> ENL3<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X13/X17/X4/M0 VREF<0> ENL3<0> VOL<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X14/X16/X3/M0 VOL<3> ENL3<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X14/X16/X4/M0 VREF<1> ENL3<1> VOL<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X14/X17/X3/M0 VOL<3> ENL3<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X14/X17/X4/M0 VREF<1> ENL3<1> VOL<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X15/X16/X3/M0 VOL<3> ENL3<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X15/X16/X4/M0 VREF<2> ENL3<2> VOL<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X15/X17/X3/M0 VOL<3> ENL3<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X120/X15/X17/X4/M0 VREF<2> ENL3<2> VOL<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X12/X14/X3/M0 X84/X121/X12/6 X84/X121/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X12/X14/X4/M0 VSS X84/X121/X12/6 X84/X121/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X12/X15/X3/M0 X84/X121/X12/7 X84/X121/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X12/X15/X4/M0 VSS X84/X121/X12/7 X84/X121/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X13/X16/X3/M0 VOL<5> ENL5<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X13/X16/X4/M0 VREF<0> ENL5<0> VOL<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X13/X17/X3/M0 VOL<5> ENL5<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X13/X17/X4/M0 VREF<0> ENL5<0> VOL<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X14/X16/X3/M0 VOL<5> ENL5<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X14/X16/X4/M0 VREF<1> ENL5<1> VOL<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X14/X17/X3/M0 VOL<5> ENL5<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X14/X17/X4/M0 VREF<1> ENL5<1> VOL<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X15/X16/X3/M0 VOL<5> ENL5<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X15/X16/X4/M0 VREF<2> ENL5<2> VOL<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X15/X17/X3/M0 VOL<5> ENL5<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X121/X15/X17/X4/M0 VREF<2> ENL5<2> VOL<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X17/X14/X3/M0 X84/X134/X17/6 X84/X134/X17/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X17/X14/X4/M0 VSS X84/X134/X17/6 X84/X134/X17/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X17/X15/X3/M0 X84/X134/X17/7 X84/X134/X17/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X17/X15/X4/M0 VSS X84/X134/X17/7 X84/X134/X17/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X24/X3/M0 VOL<6> ENL6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X24/X4/M0 VREF<0> ENL6<0> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X25/X3/M0 VOL<6> ENL6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X25/X4/M0 VREF<0> ENL6<0> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X26/X3/M0 VOL<6> ENL6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X26/X4/M0 VREF<0> ENL6<0> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X27/X3/M0 VOL<6> ENL6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X21/X27/X4/M0 VREF<0> ENL6<0> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X24/X3/M0 VOL<6> ENL6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X24/X4/M0 VREF<1> ENL6<1> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X25/X3/M0 VOL<6> ENL6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X25/X4/M0 VREF<1> ENL6<1> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X26/X3/M0 VOL<6> ENL6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X26/X4/M0 VREF<1> ENL6<1> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X27/X3/M0 VOL<6> ENL6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X22/X27/X4/M0 VREF<1> ENL6<1> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X24/X3/M0 VOL<6> ENL6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X24/X4/M0 VREF<2> ENL6<2> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X25/X3/M0 VOL<6> ENL6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X25/X4/M0 VREF<2> ENL6<2> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X26/X3/M0 VOL<6> ENL6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X26/X4/M0 VREF<2> ENL6<2> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X27/X3/M0 VOL<6> ENL6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX84/X134/X23/X27/X4/M0 VREF<2> ENL6<2> VOL<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X9/X14/X3/M0 X85/X99/X9/6 X85/X99/X9/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X9/X14/X4/M0 VSS X85/X99/X9/6 X85/X99/X9/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X9/X15/X3/M0 X85/X99/X9/7 X85/X99/X9/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X9/X15/X4/M0 VSS X85/X99/X9/7 X85/X99/X9/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X24/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X24/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X25/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X25/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X26/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X26/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X27/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X27/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X28/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X28/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X29/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X29/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X30/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X30/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X31/X3/M0 VOR<7> ENR7<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X10/X31/X4/M0 VREF<0> ENR7<0> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X24/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X24/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X25/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X25/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X26/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X26/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X27/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X27/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X28/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X28/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X29/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X29/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X30/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X30/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X31/X3/M0 VOR<7> ENR7<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X11/X31/X4/M0 VREF<1> ENR7<1> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X24/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X24/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X25/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X25/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X26/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X26/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X27/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X27/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X28/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X28/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X29/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X29/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X30/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X30/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X31/X3/M0 VOR<7> ENR7<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X99/X12/X31/X4/M0 VREF<2> ENR7<2> VOR<7> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X12/X14/X3/M0 X85/X116/X12/6 X85/X116/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X12/X14/X4/M0 VSS X85/X116/X12/6 X85/X116/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X12/X15/X3/M0 X85/X116/X12/7 X85/X116/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X12/X15/X4/M0 VSS X85/X116/X12/7 X85/X116/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X13/X16/X3/M0 VOR<0> ENR0<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X13/X16/X4/M0 VREF<0> ENR0<0> VOR<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X13/X17/X3/M0 VOR<0> ENR0<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X13/X17/X4/M0 VREF<0> ENR0<0> VOR<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X14/X16/X3/M0 VOR<0> ENR0<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X14/X16/X4/M0 VREF<1> ENR0<1> VOR<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X14/X17/X3/M0 VOR<0> ENR0<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X14/X17/X4/M0 VREF<1> ENR0<1> VOR<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X15/X16/X3/M0 VOR<0> ENR0<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X15/X16/X4/M0 VREF<2> ENR0<2> VOR<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X15/X17/X3/M0 VOR<0> ENR0<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X116/X15/X17/X4/M0 VREF<2> ENR0<2> VOR<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X12/X14/X3/M0 X85/X117/X12/6 X85/X117/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X12/X14/X4/M0 VSS X85/X117/X12/6 X85/X117/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X12/X15/X3/M0 X85/X117/X12/7 X85/X117/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X12/X15/X4/M0 VSS X85/X117/X12/7 X85/X117/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X13/X16/X3/M0 VOR<2> ENR2<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X13/X16/X4/M0 VREF<0> ENR2<0> VOR<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X13/X17/X3/M0 VOR<2> ENR2<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X13/X17/X4/M0 VREF<0> ENR2<0> VOR<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X14/X16/X3/M0 VOR<2> ENR2<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X14/X16/X4/M0 VREF<1> ENR2<1> VOR<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X14/X17/X3/M0 VOR<2> ENR2<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X14/X17/X4/M0 VREF<1> ENR2<1> VOR<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X15/X16/X3/M0 VOR<2> ENR2<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X15/X16/X4/M0 VREF<2> ENR2<2> VOR<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X15/X17/X3/M0 VOR<2> ENR2<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X117/X15/X17/X4/M0 VREF<2> ENR2<2> VOR<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X12/X14/X3/M0 X85/X118/X12/6 X85/X118/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X12/X14/X4/M0 VSS X85/X118/X12/6 X85/X118/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X12/X15/X3/M0 X85/X118/X12/7 X85/X118/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X12/X15/X4/M0 VSS X85/X118/X12/7 X85/X118/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X13/X16/X3/M0 VOR<4> ENR4<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X13/X16/X4/M0 VREF<0> ENR4<0> VOR<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X13/X17/X3/M0 VOR<4> ENR4<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X13/X17/X4/M0 VREF<0> ENR4<0> VOR<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X14/X16/X3/M0 VOR<4> ENR4<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X14/X16/X4/M0 VREF<1> ENR4<1> VOR<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X14/X17/X3/M0 VOR<4> ENR4<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X14/X17/X4/M0 VREF<1> ENR4<1> VOR<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X15/X16/X3/M0 VOR<4> ENR4<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X15/X16/X4/M0 VREF<2> ENR4<2> VOR<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X15/X17/X3/M0 VOR<4> ENR4<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X118/X15/X17/X4/M0 VREF<2> ENR4<2> VOR<4> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X12/X14/X3/M0 X85/X119/X12/6 X85/X119/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X12/X14/X4/M0 VSS X85/X119/X12/6 X85/X119/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X12/X15/X3/M0 X85/X119/X12/7 X85/X119/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X12/X15/X4/M0 VSS X85/X119/X12/7 X85/X119/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X13/X16/X3/M0 VOR<1> ENR1<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X13/X16/X4/M0 VREF<0> ENR1<0> VOR<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X13/X17/X3/M0 VOR<1> ENR1<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X13/X17/X4/M0 VREF<0> ENR1<0> VOR<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X14/X16/X3/M0 VOR<1> ENR1<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X14/X16/X4/M0 VREF<1> ENR1<1> VOR<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X14/X17/X3/M0 VOR<1> ENR1<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X14/X17/X4/M0 VREF<1> ENR1<1> VOR<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X15/X16/X3/M0 VOR<1> ENR1<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X15/X16/X4/M0 VREF<2> ENR1<2> VOR<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X15/X17/X3/M0 VOR<1> ENR1<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X119/X15/X17/X4/M0 VREF<2> ENR1<2> VOR<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X12/X14/X3/M0 X85/X120/X12/6 X85/X120/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X12/X14/X4/M0 VSS X85/X120/X12/6 X85/X120/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X12/X15/X3/M0 X85/X120/X12/7 X85/X120/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X12/X15/X4/M0 VSS X85/X120/X12/7 X85/X120/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X13/X16/X3/M0 VOR<3> ENR3<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X13/X16/X4/M0 VREF<0> ENR3<0> VOR<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X13/X17/X3/M0 VOR<3> ENR3<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X13/X17/X4/M0 VREF<0> ENR3<0> VOR<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X14/X16/X3/M0 VOR<3> ENR3<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X14/X16/X4/M0 VREF<1> ENR3<1> VOR<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X14/X17/X3/M0 VOR<3> ENR3<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X14/X17/X4/M0 VREF<1> ENR3<1> VOR<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X15/X16/X3/M0 VOR<3> ENR3<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X15/X16/X4/M0 VREF<2> ENR3<2> VOR<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X15/X17/X3/M0 VOR<3> ENR3<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X120/X15/X17/X4/M0 VREF<2> ENR3<2> VOR<3> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X12/X14/X3/M0 X85/X121/X12/6 X85/X121/X12/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X12/X14/X4/M0 VSS X85/X121/X12/6 X85/X121/X12/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X12/X15/X3/M0 X85/X121/X12/7 X85/X121/X12/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X12/X15/X4/M0 VSS X85/X121/X12/7 X85/X121/X12/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X13/X16/X3/M0 VOR<5> ENR5<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X13/X16/X4/M0 VREF<0> ENR5<0> VOR<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X13/X17/X3/M0 VOR<5> ENR5<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X13/X17/X4/M0 VREF<0> ENR5<0> VOR<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X14/X16/X3/M0 VOR<5> ENR5<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X14/X16/X4/M0 VREF<1> ENR5<1> VOR<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X14/X17/X3/M0 VOR<5> ENR5<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X14/X17/X4/M0 VREF<1> ENR5<1> VOR<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X15/X16/X3/M0 VOR<5> ENR5<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X15/X16/X4/M0 VREF<2> ENR5<2> VOR<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X15/X17/X3/M0 VOR<5> ENR5<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X121/X15/X17/X4/M0 VREF<2> ENR5<2> VOR<5> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X17/X14/X3/M0 X85/X134/X17/6 X85/X134/X17/6 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X17/X14/X4/M0 VSS X85/X134/X17/6 X85/X134/X17/6 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X17/X15/X3/M0 X85/X134/X17/7 X85/X134/X17/7 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X17/X15/X4/M0 VSS X85/X134/X17/7 X85/X134/X17/7 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X24/X3/M0 VOR<6> ENR6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X24/X4/M0 VREF<0> ENR6<0> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X25/X3/M0 VOR<6> ENR6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X25/X4/M0 VREF<0> ENR6<0> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X26/X3/M0 VOR<6> ENR6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X26/X4/M0 VREF<0> ENR6<0> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X27/X3/M0 VOR<6> ENR6<0> VREF<0> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X21/X27/X4/M0 VREF<0> ENR6<0> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X24/X3/M0 VOR<6> ENR6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X24/X4/M0 VREF<1> ENR6<1> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X25/X3/M0 VOR<6> ENR6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X25/X4/M0 VREF<1> ENR6<1> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X26/X3/M0 VOR<6> ENR6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X26/X4/M0 VREF<1> ENR6<1> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X27/X3/M0 VOR<6> ENR6<1> VREF<1> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X22/X27/X4/M0 VREF<1> ENR6<1> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X24/X3/M0 VOR<6> ENR6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X24/X4/M0 VREF<2> ENR6<2> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X25/X3/M0 VOR<6> ENR6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X25/X4/M0 VREF<2> ENR6<2> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X26/X3/M0 VOR<6> ENR6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X26/X4/M0 VREF<2> ENR6<2> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X27/X3/M0 VOR<6> ENR6<2> VREF<2> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX85/X134/X23/X27/X4/M0 VREF<2> ENR6<2> VOR<6> VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X788/X3/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X788/X4/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X789/X3/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X789/X4/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X790/X3/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X790/X4/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X791/X3/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X791/X4/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X792/X3/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X792/X4/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X793/X3/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X793/X4/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X794/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X794/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X795/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X795/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X796/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X796/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X797/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X797/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X798/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X798/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X799/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X799/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X800/X3/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X800/X4/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X801/X3/M0 X86/320 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X801/X4/M0 VSS CLKB X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X802/X3/M0 X86/320 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X802/X4/M0 VSS CLKB X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X803/X3/M0 X86/320 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X803/X4/M0 VSS CLKB X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X804/X3/M0 131 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X804/X4/M0 VSS CLKB 131 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X805/X3/M0 131 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X805/X4/M0 VSS CLKB 131 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X806/X3/M0 131 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X806/X4/M0 VSS CLKB 131 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X807/X3/M0 133 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X807/X4/M0 VSS CLKB 133 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X808/X3/M0 133 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X808/X4/M0 VSS CLKB 133 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X809/X3/M0 133 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X809/X4/M0 VSS CLKB 133 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X810/X3/M0 X86/321 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X810/X4/M0 VSS CLKB X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X811/X3/M0 X86/321 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X811/X4/M0 VSS CLKB X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X812/X3/M0 X86/321 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X812/X4/M0 VSS CLKB X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X813/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X813/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X814/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X814/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X815/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X815/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X816/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X816/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X817/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X817/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X818/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X818/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X819/X3/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X819/X4/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X820/X3/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X820/X4/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X821/X3/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X821/X4/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X822/X3/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X822/X4/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X823/X3/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X823/X4/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X824/X3/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X824/X4/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X825/X3/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X825/X4/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X971/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X971/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X972/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X972/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X973/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X973/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X974/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X974/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X975/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X975/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X976/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X976/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X977/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X977/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X978/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X978/X4/M0 131 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X979/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X979/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X980/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X980/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X981/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X981/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X982/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X982/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X983/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X983/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X984/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X984/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X985/X3/M0 VDD VDD 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X985/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X986/X3/M0 VDD VDD 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X986/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X987/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X987/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X988/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X988/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X989/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X989/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X990/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X990/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X991/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X991/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X992/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X992/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X993/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X993/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X994/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X994/X4/M0 133 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X995/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X995/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X996/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X996/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X997/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X997/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X998/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X998/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X999/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X999/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1000/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1000/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1271/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1271/X5/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1272/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1272/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1273/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1273/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1274/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1274/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1275/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1275/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1276/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1276/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1277/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1277/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1278/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1278/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1279/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1279/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1280/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1280/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1281/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1281/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1282/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1282/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1283/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1283/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1284/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1284/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1285/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1285/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1286/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1286/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1287/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1287/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1288/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1288/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1289/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1289/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1290/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1290/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1291/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1291/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1292/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1292/X5/M0 X86/325 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1293/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1293/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1294/X4/M0 131 OSP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1294/X5/M0 X86/325 OSP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1295/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1295/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1296/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1296/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1297/X4/M0 131 INP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1297/X5/M0 X86/325 INP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1298/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1298/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1299/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1299/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1300/X4/M0 131 INP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1300/X5/M0 X86/325 INP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1301/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1301/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1302/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1302/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1303/X4/M0 131 INP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1303/X5/M0 X86/325 INP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1304/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1304/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1305/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1305/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1306/X4/M0 131 INP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1306/X5/M0 X86/325 INP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1307/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1307/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1308/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1308/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1309/X4/M0 131 INP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1309/X5/M0 X86/325 INP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1310/X4/M0 X86/320 X86/321 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1310/X5/M0 131 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1311/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1311/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1312/X4/M0 131 INP X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1312/X5/M0 X86/325 INP 131 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1313/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1313/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1314/X4/M0 133 INM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1314/X5/M0 X86/325 INM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1315/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1315/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1316/X4/M0 133 INM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1316/X5/M0 X86/325 INM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1317/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1317/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1318/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1318/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1319/X4/M0 133 INM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1319/X5/M0 X86/325 INM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1320/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1320/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1321/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1321/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1322/X4/M0 133 INM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1322/X5/M0 X86/325 INM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1323/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1323/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1324/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1324/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1325/X4/M0 133 INM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1325/X5/M0 X86/325 INM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1326/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1326/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1327/X4/M0 X86/325 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1327/X5/M0 VDD CLKB X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1328/X4/M0 133 INM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1328/X5/M0 X86/325 INM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1329/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1329/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1330/X4/M0 133 OSM X86/325 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1330/X5/M0 X86/325 OSM 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1331/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1331/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1332/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1332/X5/M0 X86/325 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1333/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1333/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1334/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1334/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1335/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1335/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1336/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1336/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1337/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1337/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1338/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1338/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1339/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1339/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1340/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1340/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1341/X4/M0 X86/321 X86/320 133 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1341/X5/M0 133 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1342/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1342/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1343/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1343/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1344/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1344/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1345/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1345/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1346/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1346/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1347/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1347/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1348/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1348/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1349/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1349/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1350/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1350/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1351/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1351/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1352/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1352/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1353/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1353/X5/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1354/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1354/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
.ends


