** Schematic Netlist, pvs precompare
** 

.subckt sarafe_nsw CLKB ENL0<2> ENL0<1> ENL0<0> ENL1<2> ENL1<1> ENL1<0> ENL2<2> ENL2<1> ENL2<0> ENL3<2> ENL3<1> ENL3<0> ENL4<2> ENL4<1> ENL4<0> ENL5<2> ENL5<1> ENL5<0> ENL6<2> 
+ ENL6<1> ENL6<0> ENL7<2> ENL7<1> ENL7<0> ENR0<2> ENR0<1> ENR0<0> ENR1<2> ENR1<1> ENR1<0> ENR2<2> ENR2<1> ENR2<0> ENR3<2> ENR3<1> ENR3<0> ENR4<2> ENR4<1> ENR4<0> 
+ ENR5<2> ENR5<1> ENR5<0> ENR6<2> ENR6<1> ENR6<0> ENR7<2> ENR7<1> ENR7<0> INM INP OSM OSP OUTM OUTP VDD VOL<7> VOL<6> VOL<5> VOL<4> 
+ VOL<3> VOL<2> VOL<1> VOL<0> VOR<7> VOR<6> VOR<5> VOR<4> VOR<3> VOR<2> VOR<1> VOR<0> VREF<2> VREF<1> VREF<0> VSS 
RXICAPM0/XI7<99>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<98>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<97>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<96>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<95>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<94>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<93>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<92>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<91>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<90>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<89>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<88>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<87>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<86>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<85>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<84>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<83>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<82>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<81>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<80>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<79>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<78>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<77>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<76>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<75>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<74>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<73>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<72>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<71>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<70>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<69>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<68>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<67>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<66>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<65>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<64>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<63>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<62>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<61>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<60>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<59>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<58>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<57>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<56>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<55>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<54>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<53>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<52>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<51>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<50>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<49>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<48>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<47>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<46>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<45>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<44>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<43>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<42>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<41>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<40>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<39>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<38>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<37>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<36>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<35>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<34>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<33>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<32>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<31>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<30>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<29>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<28>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<27>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<26>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<25>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<24>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<23>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<22>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<21>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<20>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<19>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<18>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<17>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<16>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<15>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<14>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<13>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<12>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<11>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<10>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<9>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<8>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<7>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<6>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<5>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<4>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<3>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<2>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI7<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<52>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<51>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<50>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<49>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<48>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<47>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<46>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<45>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<44>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<43>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<42>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<41>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<40>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<39>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<38>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<37>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<36>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<35>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<34>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<33>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<32>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<31>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<30>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<29>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<28>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<27>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<26>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<25>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<24>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<23>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<22>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<21>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<20>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<19>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<18>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<17>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<16>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<15>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<14>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<13>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<12>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<11>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<10>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<9>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<8>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<7>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<6>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<5>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<4>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<3>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<2>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI6<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<27>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<26>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<25>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<24>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<23>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<22>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<21>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<20>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<19>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<18>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<17>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<16>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<15>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<14>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<13>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<12>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<11>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<10>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<9>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<8>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<7>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<6>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<5>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<4>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<3>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<2>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI5<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<15>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<14>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<13>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<12>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<11>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<10>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<9>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<8>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<7>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<6>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<5>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<4>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<3>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<2>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI4<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<7>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<6>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<5>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<4>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<3>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<2>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI3<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI2<3>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI2<2>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI2<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI2<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI1<1>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI1<0>/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XIC0_0/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPM0/XI0/RR0 INM INM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<99>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<98>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<97>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<96>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<95>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<94>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<93>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<92>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<91>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<90>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<89>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<88>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<87>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<86>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<85>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<84>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<83>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<82>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<81>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<80>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<79>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<78>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<77>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<76>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<75>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<74>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<73>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<72>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<71>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<70>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<69>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<68>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<67>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<66>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<65>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<64>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<63>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<62>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<61>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<60>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<59>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<58>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<57>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<56>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<55>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<54>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<53>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<52>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<51>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<50>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<49>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<48>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<47>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<46>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<45>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<44>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<43>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<42>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<41>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<40>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<39>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<38>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<37>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<36>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<35>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<34>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<33>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<32>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<31>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<30>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<29>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<28>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<27>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<26>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<25>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<24>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<23>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<22>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<21>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<20>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<19>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<18>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<17>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<16>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<15>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<14>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<13>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<12>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<11>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<10>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<9>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<8>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<7>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<6>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<5>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<4>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<3>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<2>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI7<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<52>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<51>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<50>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<49>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<48>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<47>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<46>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<45>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<44>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<43>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<42>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<41>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<40>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<39>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<38>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<37>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<36>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<35>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<34>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<33>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<32>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<31>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<30>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<29>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<28>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<27>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<26>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<25>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<24>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<23>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<22>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<21>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<20>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<19>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<18>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<17>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<16>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<15>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<14>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<13>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<12>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<11>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<10>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<9>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<8>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<7>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<6>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<5>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<4>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<3>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<2>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI6<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<27>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<26>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<25>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<24>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<23>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<22>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<21>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<20>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<19>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<18>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<17>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<16>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<15>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<14>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<13>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<12>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<11>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<10>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<9>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<8>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<7>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<6>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<5>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<4>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<3>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<2>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI5<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<15>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<14>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<13>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<12>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<11>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<10>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<9>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<8>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<7>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<6>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<5>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<4>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<3>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<2>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI4<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<7>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<6>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<5>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<4>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<3>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<2>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI3<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI2<3>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI2<2>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI2<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI2<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI1<1>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI1<0>/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XIC0_0/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXICAPP0/XI0/RR0 INP INP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
MXISA0/XIRGNNDM1/MM0 XISA0/OP XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIBUFN0/MM0 OUTP XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIBUFN1/MM0 OUTM XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIRST1/MM0 INTP CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRST3/MM0 XISA0/OP CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRST0/MM0 INTM CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRST2/MM0 XISA0/OM CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRGNNDM0/MM0 XISA0/OM XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIRGNN0/MM0 XISA0/OM XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIRGNN1/MM0 XISA0/OP XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIBUFP0/MM0 OUTP XISA0/OM VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIBUFP1/MM0 OUTM XISA0/OP VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIRGNPDM2/MM0 INTP VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIRGNPDM1/MM0 INTM VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIRGNPDM0/MM0 VDD VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISA0/XIRGNP1/MM0 XISA0/OP XISA0/OM INTP VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=22 
MXISA0/XIRGNP0/MM0 XISA0/OM XISA0/OP INTM VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=22 
MXISA0/XIOSM0/MM0 INTP OSM XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIOSP0/MM0 INTM OSP XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIOSPB0/MM0 VDD OSP VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=20 
MXISA0/XIOSMB0/MM0 VDD OSM VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=20 
MXISA0/XIINDM1/MM0 VDD VDD XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIINDM0/MM0 VDD VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XICKPDM0/MM0 VDD VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=52 
MXISA0/XICKP0/MM0 XISA0/TAIL CLKB VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=24 
MXISA0/XIINM0/MM0 INTP INM XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIINP0/MM0 INTM INP XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXICDRVM0/XICDRV3/XISW0/XIN1/MM0 VREF<2> ENR3<2> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW0/XIN0/MM0 VREF<2> ENR3<2> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW1/XIN1/MM0 VREF<1> ENR3<1> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW1/XIN0/MM0 VREF<1> ENR3<1> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW2/XIN1/MM0 VREF<0> ENR3<0> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW2/XIN0/MM0 VREF<0> ENR3<0> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XITIE0/XIN1/MM0 XICDRVM0/XICDRV3/XITIE0/net5 XICDRVM0/XICDRV3/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XITIE0/XIN0/MM0 XICDRVM0/XICDRV3/XITIE0/net6 XICDRVM0/XICDRV3/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW0/XIN1/MM0 VREF<2> ENR0<2> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW0/XIN0/MM0 VREF<2> ENR0<2> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW1/XIN1/MM0 VREF<1> ENR0<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW1/XIN0/MM0 VREF<1> ENR0<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW2/XIN1/MM0 VREF<0> ENR0<0> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW2/XIN0/MM0 VREF<0> ENR0<0> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XITIE0/XIN1/MM0 XICDRVM0/XICDRV0/XITIE0/net5 XICDRVM0/XICDRV0/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XITIE0/XIN0/MM0 XICDRVM0/XICDRV0/XITIE0/net6 XICDRVM0/XICDRV0/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW0/XIN1/MM0 VREF<2> ENR2<2> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW0/XIN0/MM0 VREF<2> ENR2<2> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW1/XIN1/MM0 VREF<1> ENR2<1> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW1/XIN0/MM0 VREF<1> ENR2<1> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW2/XIN1/MM0 VREF<0> ENR2<0> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW2/XIN0/MM0 VREF<0> ENR2<0> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XITIE0/XIN1/MM0 XICDRVM0/XICDRV2/XITIE0/net5 XICDRVM0/XICDRV2/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XITIE0/XIN0/MM0 XICDRVM0/XICDRV2/XITIE0/net6 XICDRVM0/XICDRV2/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW0/XIN1/MM0 VREF<2> ENR1<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW0/XIN0/MM0 VREF<2> ENR1<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW1/XIN1/MM0 VREF<1> ENR1<1> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW1/XIN0/MM0 VREF<1> ENR1<1> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW2/XIN1/MM0 VREF<0> ENR1<0> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW2/XIN0/MM0 VREF<0> ENR1<0> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XITIE0/XIN1/MM0 XICDRVM0/XICDRV1/XITIE0/net5 XICDRVM0/XICDRV1/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XITIE0/XIN0/MM0 XICDRVM0/XICDRV1/XITIE0/net6 XICDRVM0/XICDRV1/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW0/XIN1/MM0 VREF<2> ENR4<2> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW0/XIN0/MM0 VREF<2> ENR4<2> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW1/XIN1/MM0 VREF<1> ENR4<1> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW1/XIN0/MM0 VREF<1> ENR4<1> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW2/XIN1/MM0 VREF<0> ENR4<0> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW2/XIN0/MM0 VREF<0> ENR4<0> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XITIE0/XIN1/MM0 XICDRVM0/XICDRV4/XITIE0/net5 XICDRVM0/XICDRV4/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XITIE0/XIN0/MM0 XICDRVM0/XICDRV4/XITIE0/net6 XICDRVM0/XICDRV4/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW0/XIN1/MM0 VREF<2> ENR5<2> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW0/XIN0/MM0 VREF<2> ENR5<2> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW1/XIN1/MM0 VREF<1> ENR5<1> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW1/XIN0/MM0 VREF<1> ENR5<1> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW2/XIN1/MM0 VREF<0> ENR5<0> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW2/XIN0/MM0 VREF<0> ENR5<0> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XITIE0/XIN1/MM0 XICDRVM0/XICDRV5/XITIE0/net5 XICDRVM0/XICDRV5/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XITIE0/XIN0/MM0 XICDRVM0/XICDRV5/XITIE0/net6 XICDRVM0/XICDRV5/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV6/XITIE0/XIN1/MM0 XICDRVM0/XICDRV6/XITIE0/net5 XICDRVM0/XICDRV6/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV6/XITIE0/XIN0/MM0 XICDRVM0/XICDRV6/XITIE0/net6 XICDRVM0/XICDRV6/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV6/XISW0/XIN1/MM0 VREF<2> ENR6<2> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW0/XIN0/MM0 VREF<2> ENR6<2> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW1/XIN1/MM0 VREF<1> ENR6<1> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW1/XIN0/MM0 VREF<1> ENR6<1> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW2/XIN1/MM0 VREF<0> ENR6<0> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW2/XIN0/MM0 VREF<0> ENR6<0> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV7/XITIE0/XIN1/MM0 XICDRVM0/XICDRV7/XITIE0/net5 XICDRVM0/XICDRV7/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV7/XITIE0/XIN0/MM0 XICDRVM0/XICDRV7/XITIE0/net6 XICDRVM0/XICDRV7/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV7/XISW0/XIN1/MM0 VREF<2> ENR7<2> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW0/XIN0/MM0 VREF<2> ENR7<2> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW1/XIN1/MM0 VREF<1> ENR7<1> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW1/XIN0/MM0 VREF<1> ENR7<1> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW2/XIN1/MM0 VREF<0> ENR7<0> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW2/XIN0/MM0 VREF<0> ENR7<0> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV3/XISW0/XIN1/MM0 VREF<2> ENL3<2> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW0/XIN0/MM0 VREF<2> ENL3<2> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW1/XIN1/MM0 VREF<1> ENL3<1> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW1/XIN0/MM0 VREF<1> ENL3<1> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW2/XIN1/MM0 VREF<0> ENL3<0> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW2/XIN0/MM0 VREF<0> ENL3<0> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XITIE0/XIN1/MM0 XICDRVP0/XICDRV3/XITIE0/net5 XICDRVP0/XICDRV3/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XITIE0/XIN0/MM0 XICDRVP0/XICDRV3/XITIE0/net6 XICDRVP0/XICDRV3/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW0/XIN1/MM0 VREF<2> ENL0<2> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW0/XIN0/MM0 VREF<2> ENL0<2> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW1/XIN1/MM0 VREF<1> ENL0<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW1/XIN0/MM0 VREF<1> ENL0<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW2/XIN1/MM0 VREF<0> ENL0<0> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW2/XIN0/MM0 VREF<0> ENL0<0> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XITIE0/XIN1/MM0 XICDRVP0/XICDRV0/XITIE0/net5 XICDRVP0/XICDRV0/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XITIE0/XIN0/MM0 XICDRVP0/XICDRV0/XITIE0/net6 XICDRVP0/XICDRV0/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW0/XIN1/MM0 VREF<2> ENL2<2> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW0/XIN0/MM0 VREF<2> ENL2<2> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW1/XIN1/MM0 VREF<1> ENL2<1> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW1/XIN0/MM0 VREF<1> ENL2<1> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW2/XIN1/MM0 VREF<0> ENL2<0> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW2/XIN0/MM0 VREF<0> ENL2<0> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XITIE0/XIN1/MM0 XICDRVP0/XICDRV2/XITIE0/net5 XICDRVP0/XICDRV2/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XITIE0/XIN0/MM0 XICDRVP0/XICDRV2/XITIE0/net6 XICDRVP0/XICDRV2/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW0/XIN1/MM0 VREF<2> ENL1<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW0/XIN0/MM0 VREF<2> ENL1<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW1/XIN1/MM0 VREF<1> ENL1<1> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW1/XIN0/MM0 VREF<1> ENL1<1> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW2/XIN1/MM0 VREF<0> ENL1<0> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW2/XIN0/MM0 VREF<0> ENL1<0> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XITIE0/XIN1/MM0 XICDRVP0/XICDRV1/XITIE0/net5 XICDRVP0/XICDRV1/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XITIE0/XIN0/MM0 XICDRVP0/XICDRV1/XITIE0/net6 XICDRVP0/XICDRV1/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW0/XIN1/MM0 VREF<2> ENL4<2> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW0/XIN0/MM0 VREF<2> ENL4<2> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW1/XIN1/MM0 VREF<1> ENL4<1> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW1/XIN0/MM0 VREF<1> ENL4<1> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW2/XIN1/MM0 VREF<0> ENL4<0> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW2/XIN0/MM0 VREF<0> ENL4<0> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XITIE0/XIN1/MM0 XICDRVP0/XICDRV4/XITIE0/net5 XICDRVP0/XICDRV4/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XITIE0/XIN0/MM0 XICDRVP0/XICDRV4/XITIE0/net6 XICDRVP0/XICDRV4/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW0/XIN1/MM0 VREF<2> ENL5<2> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW0/XIN0/MM0 VREF<2> ENL5<2> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW1/XIN1/MM0 VREF<1> ENL5<1> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW1/XIN0/MM0 VREF<1> ENL5<1> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW2/XIN1/MM0 VREF<0> ENL5<0> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW2/XIN0/MM0 VREF<0> ENL5<0> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XITIE0/XIN1/MM0 XICDRVP0/XICDRV5/XITIE0/net5 XICDRVP0/XICDRV5/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XITIE0/XIN0/MM0 XICDRVP0/XICDRV5/XITIE0/net6 XICDRVP0/XICDRV5/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV6/XITIE0/XIN1/MM0 XICDRVP0/XICDRV6/XITIE0/net5 XICDRVP0/XICDRV6/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV6/XITIE0/XIN0/MM0 XICDRVP0/XICDRV6/XITIE0/net6 XICDRVP0/XICDRV6/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV6/XISW0/XIN1/MM0 VREF<2> ENL6<2> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW0/XIN0/MM0 VREF<2> ENL6<2> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW1/XIN1/MM0 VREF<1> ENL6<1> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW1/XIN0/MM0 VREF<1> ENL6<1> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW2/XIN1/MM0 VREF<0> ENL6<0> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW2/XIN0/MM0 VREF<0> ENL6<0> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV7/XITIE0/XIN1/MM0 XICDRVP0/XICDRV7/XITIE0/net5 XICDRVP0/XICDRV7/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV7/XITIE0/XIN0/MM0 XICDRVP0/XICDRV7/XITIE0/net6 XICDRVP0/XICDRV7/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV7/XISW0/XIN1/MM0 VREF<2> ENL7<2> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW0/XIN0/MM0 VREF<2> ENL7<2> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW1/XIN1/MM0 VREF<1> ENL7<1> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW1/XIN0/MM0 VREF<1> ENL7<1> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW2/XIN1/MM0 VREF<0> ENL7<0> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW2/XIN0/MM0 VREF<0> ENL7<0> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
.ends


