** Layout Netlist, pvs precompare
** 

.subckt sarafe_nsw CLKB ENL0<0> ENL0<1> ENL0<2> ENL1<0> ENL1<1> ENL1<2> ENL2<0> ENL2<1> ENL2<2> ENL3<0> ENL3<1> ENL3<2> ENL4<0> ENL4<1> ENL4<2> ENL5<0> ENL5<1> ENL5<2> ENL6<0> 
+ ENL6<1> ENL6<2> ENL7<0> ENL7<1> ENL7<2> ENR0<0> ENR0<1> ENR0<2> ENR1<0> ENR1<1> ENR1<2> ENR2<0> ENR2<1> ENR2<2> ENR3<0> ENR3<1> ENR3<2> ENR4<0> ENR4<1> ENR4<2> 
+ ENR5<0> ENR5<1> ENR5<2> ENR6<0> ENR6<1> ENR6<2> ENR7<0> ENR7<1> ENR7<2> INM INP OSM OSP OUTM OUTP VDD VOL<0> VOL<1> VOL<2> VOL<3> 
+ VOL<4> VOL<5> VOL<6> VOL<7> VOR<0> VOR<1> VOR<2> VOR<3> VOR<4> VOR<5> VOR<6> VOR<7> VREF<0> VREF<1> VREF<2> VSS 
RX82/X50/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X51/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X52/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X53/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X54/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X55/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X56/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X57/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X58/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X59/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X60/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X61/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X62/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X63/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X64/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X65/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X66/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X67/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X68/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X69/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X70/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X71/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X72/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X73/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X74/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X75/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X76/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X77/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X78/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X79/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X80/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X81/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X82/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X83/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X84/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X85/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X86/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X87/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X88/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X89/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X90/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X91/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X92/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X93/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X94/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X95/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X96/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X97/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X98/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X99/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X100/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X101/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X102/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X103/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X104/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X105/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X106/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X107/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X108/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X109/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X110/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X111/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X112/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X113/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X114/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X115/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X116/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X117/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X118/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X119/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X120/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X121/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X122/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X123/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X124/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X125/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X126/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X127/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X128/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X129/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X130/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X131/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X132/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X133/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X134/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X135/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X136/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X137/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X138/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X139/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X140/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X141/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X142/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X143/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X144/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X145/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X146/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X147/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X148/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X149/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X150/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X151/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X152/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X153/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X154/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X155/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X156/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X157/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X158/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X159/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X160/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X161/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X162/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X163/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X164/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X165/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X166/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X167/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X168/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X169/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X170/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X171/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X172/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X173/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X174/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X175/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X176/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X177/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X178/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X179/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X180/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X181/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X182/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X183/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X184/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X185/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X186/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X187/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X188/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X189/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X190/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X191/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X192/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X193/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X194/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X195/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X196/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X197/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X198/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X199/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X200/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X201/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X202/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X203/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X204/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X205/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X206/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X207/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X208/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X209/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X210/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X211/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X212/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X213/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X214/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X215/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X216/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X217/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X218/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X219/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X220/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X221/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X222/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X223/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X224/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X225/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X226/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X227/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X228/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X229/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X230/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X231/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X232/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X233/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X234/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X235/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X236/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X237/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X238/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X239/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X240/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X241/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X242/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X243/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X244/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X245/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X246/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X247/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X248/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X249/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X250/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X251/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X252/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X253/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X254/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X255/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X256/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X257/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X258/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X259/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X260/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X261/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX82/X262/R0 INP INP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X50/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X51/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X52/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X53/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X54/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X55/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X56/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X57/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X58/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X59/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X60/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X61/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X62/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X63/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X64/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X65/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X66/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X67/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X68/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X69/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X70/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X71/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X72/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X73/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X74/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X75/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X76/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X77/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X78/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X79/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X80/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X81/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X82/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X83/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X84/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X85/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X86/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X87/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X88/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X89/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X90/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X91/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X92/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X93/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X94/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X95/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X96/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X97/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X98/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X99/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X100/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X101/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X102/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X103/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X104/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X105/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X106/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X107/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X108/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X109/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X110/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X111/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X112/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X113/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X114/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X115/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X116/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X117/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X118/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X119/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X120/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X121/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X122/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X123/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X124/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X125/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X126/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X127/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X128/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X129/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X130/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X131/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X132/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X133/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X134/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X135/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X136/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X137/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X138/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X139/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X140/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X141/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X142/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X143/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X144/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X145/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X146/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X147/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X148/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X149/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X150/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X151/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X152/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X153/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X154/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X155/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X156/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X157/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X158/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X159/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X160/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X161/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X162/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X163/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X164/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X165/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X166/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X167/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X168/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X169/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X170/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X171/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X172/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X173/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X174/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X175/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X176/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X177/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X178/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X179/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X180/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X181/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X182/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X183/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X184/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X185/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X186/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X187/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X188/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X189/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X190/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X191/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X192/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X193/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X194/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X195/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X196/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X197/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X198/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X199/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X200/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X201/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X202/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X203/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X204/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X205/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X206/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X207/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X208/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X209/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X210/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X211/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X212/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X213/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X214/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X215/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X216/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X217/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X218/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X219/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X220/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X221/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X222/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X223/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X224/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X225/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X226/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X227/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X228/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X229/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X230/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X231/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X232/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X233/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X234/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X235/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X236/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X237/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X238/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X239/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X240/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X241/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X242/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X243/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X244/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X245/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X246/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X247/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X248/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X249/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X250/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X251/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X252/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X253/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X254/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X255/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X256/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X257/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X258/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X259/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X260/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X261/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX83/X262/R0 INM INM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
MX86/X791/X0/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X791/X1/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X792/X0/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X792/X1/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X793/X0/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X793/X1/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X794/X0/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X794/X1/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X795/X0/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X795/X1/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X796/X0/M0 OUTP X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X796/X1/M0 VSS X86/320 OUTP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X797/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X797/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X798/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X798/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X799/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X799/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X800/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X800/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X801/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X801/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X802/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X802/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X803/X0/M0 X86/320 X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X803/X1/M0 VSS X86/321 X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X804/X0/M0 X86/320 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X804/X1/M0 VSS CLKB X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X805/X0/M0 X86/320 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X805/X1/M0 VSS CLKB X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X806/X0/M0 X86/320 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X806/X1/M0 VSS CLKB X86/320 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X807/X0/M0 87 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X807/X1/M0 VSS CLKB 87 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X808/X0/M0 87 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X808/X1/M0 VSS CLKB 87 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X809/X0/M0 87 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X809/X1/M0 VSS CLKB 87 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X810/X0/M0 89 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X810/X1/M0 VSS CLKB 89 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X811/X0/M0 89 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X811/X1/M0 VSS CLKB 89 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X812/X0/M0 89 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X812/X1/M0 VSS CLKB 89 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X813/X0/M0 X86/321 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X813/X1/M0 VSS CLKB X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X814/X0/M0 X86/321 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X814/X1/M0 VSS CLKB X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X815/X0/M0 X86/321 CLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X815/X1/M0 VSS CLKB X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X816/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X816/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X817/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X817/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X818/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X818/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X819/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X819/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X820/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X820/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X821/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X821/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X822/X0/M0 X86/321 X86/320 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X822/X1/M0 VSS X86/320 X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X823/X0/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X823/X1/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X824/X0/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X824/X1/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X825/X0/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X825/X1/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X826/X0/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X826/X1/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X827/X0/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X827/X1/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X828/X0/M0 OUTM X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X828/X1/M0 VSS X86/321 OUTM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X941/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X941/X5/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X942/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X942/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X943/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X943/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X944/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X944/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X945/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X945/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X946/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X946/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X947/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X947/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X948/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X948/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X949/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X949/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X950/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X950/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X951/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X951/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X952/X4/M0 OUTP X86/320 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X952/X5/M0 VDD X86/320 OUTP VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X953/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X953/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X954/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X954/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X955/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X955/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X956/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X956/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X957/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X957/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X958/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X958/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X959/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X959/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X960/X4/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X960/X5/M0 VDD OSP VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X961/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X961/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X962/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X962/X5/M0 X86/324 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X963/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X963/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X964/X4/M0 87 OSP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X964/X5/M0 X86/324 OSP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X965/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X965/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X966/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X966/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X967/X4/M0 87 INP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X967/X5/M0 X86/324 INP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X968/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X968/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X969/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X969/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X970/X4/M0 87 INP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X970/X5/M0 X86/324 INP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X971/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X971/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X972/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X972/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X973/X4/M0 87 INP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X973/X5/M0 X86/324 INP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X974/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X974/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X975/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X975/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X976/X4/M0 87 INP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X976/X5/M0 X86/324 INP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X977/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X977/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X978/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X978/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X979/X4/M0 87 INP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X979/X5/M0 X86/324 INP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X980/X4/M0 X86/320 X86/321 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X980/X5/M0 87 X86/321 X86/320 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X981/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X981/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X982/X4/M0 87 INP X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X982/X5/M0 X86/324 INP 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X983/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X983/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X984/X4/M0 89 INM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X984/X5/M0 X86/324 INM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X985/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X985/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X986/X4/M0 89 INM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X986/X5/M0 X86/324 INM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X987/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X987/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X988/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X988/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X989/X4/M0 89 INM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X989/X5/M0 X86/324 INM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X990/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X990/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X991/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X991/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X992/X4/M0 89 INM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X992/X5/M0 X86/324 INM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X993/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X993/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X994/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X994/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X995/X4/M0 89 INM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X995/X5/M0 X86/324 INM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X996/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X996/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X997/X4/M0 X86/324 CLKB VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X997/X5/M0 VDD CLKB X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X998/X4/M0 89 INM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X998/X5/M0 X86/324 INM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X999/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X999/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1000/X4/M0 89 OSM X86/324 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1000/X5/M0 X86/324 OSM 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1001/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1001/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1002/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1002/X5/M0 X86/324 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1003/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1003/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1004/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1004/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1005/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1005/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1006/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1006/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1007/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1007/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1008/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1008/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1009/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1009/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1010/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1010/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1011/X4/M0 X86/321 X86/320 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1011/X5/M0 89 X86/320 X86/321 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1012/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1012/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1013/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1013/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1014/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1014/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1015/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1015/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1016/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1016/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1017/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1017/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1018/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1018/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1019/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1019/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1020/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1020/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1021/X4/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1021/X5/M0 VDD OSM VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1022/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1022/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1023/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1023/X5/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1024/X4/M0 OUTM X86/321 VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1024/X5/M0 VDD X86/321 OUTM VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1390/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1390/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1391/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1391/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1392/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1392/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1393/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1393/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1394/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1394/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1395/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1395/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1396/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1396/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1397/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1397/X4/M0 87 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1398/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1398/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1399/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1399/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1400/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1400/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1401/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1401/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1402/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1402/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1403/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1403/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1404/X3/M0 VDD VDD 87 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1404/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1405/X3/M0 VDD VDD 89 VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1405/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1406/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1406/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1407/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1407/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1408/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1408/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1409/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1409/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1410/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1410/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1411/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1411/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1412/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1412/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1413/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1413/X4/M0 89 VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1414/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1414/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1415/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1415/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1416/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1416/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1417/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1417/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1418/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1418/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1419/X3/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX86/X1419/X4/M0 VDD VDD VDD VDD P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
.ends


