** Schematic Netlist, pvs precompare
** 

.subckt sarafe_nsw CLKB ENL0<2> ENL0<1> ENL0<0> ENL1<2> ENL1<1> ENL1<0> ENL2<2> ENL2<1> ENL2<0> ENL3<2> ENL3<1> ENL3<0> ENL4<2> ENL4<1> ENL4<0> ENL5<2> ENL5<1> ENL5<0> ENL6<2> 
+ ENL6<1> ENL6<0> ENL7<2> ENL7<1> ENL7<0> ENR0<2> ENR0<1> ENR0<0> ENR1<2> ENR1<1> ENR1<0> ENR2<2> ENR2<1> ENR2<0> ENR3<2> ENR3<1> ENR3<0> ENR4<2> ENR4<1> ENR4<0> 
+ ENR5<2> ENR5<1> ENR5<0> ENR6<2> ENR6<1> ENR6<0> ENR7<2> ENR7<1> ENR7<0> INM INP OSM OSP OUTM OUTP VDD VOL<7> VOL<6> VOL<5> VOL<4> 
+ VOL<3> VOL<2> VOL<1> VOL<0> VOR<7> VOR<6> VOR<5> VOR<4> VOR<3> VOR<2> VOR<1> VOR<0> VREF<2> VREF<1> VREF<0> VSS 
MXISA0/XIRGNNDM1/MM0 XISA0/OP XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIBUFN0/MM0 OUTP XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIBUFN1/MM0 OUTM XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIRST1/MM0 INTP CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRST3/MM0 XISA0/OP CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRST0/MM0 INTM CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRST2/MM0 XISA0/OM CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XIRGNNDM0/MM0 XISA0/OM XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIRGNN0/MM0 XISA0/OM XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIRGNN1/MM0 XISA0/OP XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIBUFP0/MM0 OUTP XISA0/OM VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIBUFP1/MM0 OUTM XISA0/OP VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIRGNPDM2/MM0 INTP VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIRGNPDM1/MM0 INTM VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIRGNPDM0/MM0 VDD VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISA0/XIRGNP1/MM0 XISA0/OP XISA0/OM INTP VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=22 
MXISA0/XIRGNP0/MM0 XISA0/OM XISA0/OP INTM VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=22 
MXISA0/XIOSM0/MM0 INTP OSM XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIOSP0/MM0 INTM OSP XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIOSPB0/MM0 VDD OSP VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=20 
MXISA0/XIOSMB0/MM0 VDD OSM VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=20 
MXISA0/XIINDM1/MM0 VDD VDD XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISA0/XIINDM0/MM0 VDD VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISA0/XICKPDM0/MM0 VDD VDD VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=52 
MXISA0/XICKP0/MM0 XISA0/TAIL CLKB VDD VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=24 
MXISA0/XIINM0/MM0 INTP INM XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISA0/XIINP0/MM0 INTM INP XISA0/TAIL VDD P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXICDRVM0/XICDRV3/XISW0/XIN1/MM0 VREF<2> ENR3<2> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW0/XIN0/MM0 VREF<2> ENR3<2> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW1/XIN1/MM0 VREF<1> ENR3<1> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW1/XIN0/MM0 VREF<1> ENR3<1> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW2/XIN1/MM0 VREF<0> ENR3<0> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XISW2/XIN0/MM0 VREF<0> ENR3<0> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XITIE0/XIN1/MM0 XICDRVM0/XICDRV3/XITIE0/net5 XICDRVM0/XICDRV3/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV3/XITIE0/XIN0/MM0 XICDRVM0/XICDRV3/XITIE0/net6 XICDRVM0/XICDRV3/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW0/XIN1/MM0 VREF<2> ENR0<2> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW0/XIN0/MM0 VREF<2> ENR0<2> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW1/XIN1/MM0 VREF<1> ENR0<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW1/XIN0/MM0 VREF<1> ENR0<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW2/XIN1/MM0 VREF<0> ENR0<0> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XISW2/XIN0/MM0 VREF<0> ENR0<0> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XITIE0/XIN1/MM0 XICDRVM0/XICDRV0/XITIE0/net5 XICDRVM0/XICDRV0/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV0/XITIE0/XIN0/MM0 XICDRVM0/XICDRV0/XITIE0/net6 XICDRVM0/XICDRV0/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW0/XIN1/MM0 VREF<2> ENR2<2> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW0/XIN0/MM0 VREF<2> ENR2<2> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW1/XIN1/MM0 VREF<1> ENR2<1> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW1/XIN0/MM0 VREF<1> ENR2<1> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW2/XIN1/MM0 VREF<0> ENR2<0> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XISW2/XIN0/MM0 VREF<0> ENR2<0> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XITIE0/XIN1/MM0 XICDRVM0/XICDRV2/XITIE0/net5 XICDRVM0/XICDRV2/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV2/XITIE0/XIN0/MM0 XICDRVM0/XICDRV2/XITIE0/net6 XICDRVM0/XICDRV2/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW0/XIN1/MM0 VREF<2> ENR1<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW0/XIN0/MM0 VREF<2> ENR1<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW1/XIN1/MM0 VREF<1> ENR1<1> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW1/XIN0/MM0 VREF<1> ENR1<1> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW2/XIN1/MM0 VREF<0> ENR1<0> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XISW2/XIN0/MM0 VREF<0> ENR1<0> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XITIE0/XIN1/MM0 XICDRVM0/XICDRV1/XITIE0/net5 XICDRVM0/XICDRV1/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV1/XITIE0/XIN0/MM0 XICDRVM0/XICDRV1/XITIE0/net6 XICDRVM0/XICDRV1/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW0/XIN1/MM0 VREF<2> ENR4<2> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW0/XIN0/MM0 VREF<2> ENR4<2> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW1/XIN1/MM0 VREF<1> ENR4<1> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW1/XIN0/MM0 VREF<1> ENR4<1> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW2/XIN1/MM0 VREF<0> ENR4<0> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XISW2/XIN0/MM0 VREF<0> ENR4<0> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XITIE0/XIN1/MM0 XICDRVM0/XICDRV4/XITIE0/net5 XICDRVM0/XICDRV4/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV4/XITIE0/XIN0/MM0 XICDRVM0/XICDRV4/XITIE0/net6 XICDRVM0/XICDRV4/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW0/XIN1/MM0 VREF<2> ENR5<2> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW0/XIN0/MM0 VREF<2> ENR5<2> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW1/XIN1/MM0 VREF<1> ENR5<1> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW1/XIN0/MM0 VREF<1> ENR5<1> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW2/XIN1/MM0 VREF<0> ENR5<0> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XISW2/XIN0/MM0 VREF<0> ENR5<0> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XITIE0/XIN1/MM0 XICDRVM0/XICDRV5/XITIE0/net5 XICDRVM0/XICDRV5/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV5/XITIE0/XIN0/MM0 XICDRVM0/XICDRV5/XITIE0/net6 XICDRVM0/XICDRV5/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV6/XITIE0/XIN1/MM0 XICDRVM0/XICDRV6/XITIE0/net5 XICDRVM0/XICDRV6/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV6/XITIE0/XIN0/MM0 XICDRVM0/XICDRV6/XITIE0/net6 XICDRVM0/XICDRV6/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV6/XISW0/XIN1/MM0 VREF<2> ENR6<2> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW0/XIN0/MM0 VREF<2> ENR6<2> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW1/XIN1/MM0 VREF<1> ENR6<1> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW1/XIN0/MM0 VREF<1> ENR6<1> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW2/XIN1/MM0 VREF<0> ENR6<0> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV6/XISW2/XIN0/MM0 VREF<0> ENR6<0> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVM0/XICDRV7/XITIE0/XIN1/MM0 XICDRVM0/XICDRV7/XITIE0/net5 XICDRVM0/XICDRV7/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV7/XITIE0/XIN0/MM0 XICDRVM0/XICDRV7/XITIE0/net6 XICDRVM0/XICDRV7/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVM0/XICDRV7/XISW0/XIN1/MM0 VREF<2> ENR7<2> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW0/XIN0/MM0 VREF<2> ENR7<2> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW1/XIN1/MM0 VREF<1> ENR7<1> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW1/XIN0/MM0 VREF<1> ENR7<1> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW2/XIN1/MM0 VREF<0> ENR7<0> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVM0/XICDRV7/XISW2/XIN0/MM0 VREF<0> ENR7<0> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV3/XISW0/XIN1/MM0 VREF<2> ENL3<2> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW0/XIN0/MM0 VREF<2> ENL3<2> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW1/XIN1/MM0 VREF<1> ENL3<1> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW1/XIN0/MM0 VREF<1> ENL3<1> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW2/XIN1/MM0 VREF<0> ENL3<0> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XISW2/XIN0/MM0 VREF<0> ENL3<0> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XITIE0/XIN1/MM0 XICDRVP0/XICDRV3/XITIE0/net5 XICDRVP0/XICDRV3/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV3/XITIE0/XIN0/MM0 XICDRVP0/XICDRV3/XITIE0/net6 XICDRVP0/XICDRV3/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW0/XIN1/MM0 VREF<2> ENL0<2> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW0/XIN0/MM0 VREF<2> ENL0<2> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW1/XIN1/MM0 VREF<1> ENL0<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW1/XIN0/MM0 VREF<1> ENL0<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW2/XIN1/MM0 VREF<0> ENL0<0> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XISW2/XIN0/MM0 VREF<0> ENL0<0> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XITIE0/XIN1/MM0 XICDRVP0/XICDRV0/XITIE0/net5 XICDRVP0/XICDRV0/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV0/XITIE0/XIN0/MM0 XICDRVP0/XICDRV0/XITIE0/net6 XICDRVP0/XICDRV0/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW0/XIN1/MM0 VREF<2> ENL2<2> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW0/XIN0/MM0 VREF<2> ENL2<2> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW1/XIN1/MM0 VREF<1> ENL2<1> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW1/XIN0/MM0 VREF<1> ENL2<1> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW2/XIN1/MM0 VREF<0> ENL2<0> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XISW2/XIN0/MM0 VREF<0> ENL2<0> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XITIE0/XIN1/MM0 XICDRVP0/XICDRV2/XITIE0/net5 XICDRVP0/XICDRV2/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV2/XITIE0/XIN0/MM0 XICDRVP0/XICDRV2/XITIE0/net6 XICDRVP0/XICDRV2/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW0/XIN1/MM0 VREF<2> ENL1<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW0/XIN0/MM0 VREF<2> ENL1<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW1/XIN1/MM0 VREF<1> ENL1<1> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW1/XIN0/MM0 VREF<1> ENL1<1> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW2/XIN1/MM0 VREF<0> ENL1<0> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XISW2/XIN0/MM0 VREF<0> ENL1<0> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XITIE0/XIN1/MM0 XICDRVP0/XICDRV1/XITIE0/net5 XICDRVP0/XICDRV1/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV1/XITIE0/XIN0/MM0 XICDRVP0/XICDRV1/XITIE0/net6 XICDRVP0/XICDRV1/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW0/XIN1/MM0 VREF<2> ENL4<2> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW0/XIN0/MM0 VREF<2> ENL4<2> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW1/XIN1/MM0 VREF<1> ENL4<1> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW1/XIN0/MM0 VREF<1> ENL4<1> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW2/XIN1/MM0 VREF<0> ENL4<0> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XISW2/XIN0/MM0 VREF<0> ENL4<0> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XITIE0/XIN1/MM0 XICDRVP0/XICDRV4/XITIE0/net5 XICDRVP0/XICDRV4/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV4/XITIE0/XIN0/MM0 XICDRVP0/XICDRV4/XITIE0/net6 XICDRVP0/XICDRV4/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW0/XIN1/MM0 VREF<2> ENL5<2> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW0/XIN0/MM0 VREF<2> ENL5<2> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW1/XIN1/MM0 VREF<1> ENL5<1> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW1/XIN0/MM0 VREF<1> ENL5<1> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW2/XIN1/MM0 VREF<0> ENL5<0> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XISW2/XIN0/MM0 VREF<0> ENL5<0> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XITIE0/XIN1/MM0 XICDRVP0/XICDRV5/XITIE0/net5 XICDRVP0/XICDRV5/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV5/XITIE0/XIN0/MM0 XICDRVP0/XICDRV5/XITIE0/net6 XICDRVP0/XICDRV5/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV6/XITIE0/XIN1/MM0 XICDRVP0/XICDRV6/XITIE0/net5 XICDRVP0/XICDRV6/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV6/XITIE0/XIN0/MM0 XICDRVP0/XICDRV6/XITIE0/net6 XICDRVP0/XICDRV6/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV6/XISW0/XIN1/MM0 VREF<2> ENL6<2> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW0/XIN0/MM0 VREF<2> ENL6<2> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW1/XIN1/MM0 VREF<1> ENL6<1> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW1/XIN0/MM0 VREF<1> ENL6<1> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW2/XIN1/MM0 VREF<0> ENL6<0> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV6/XISW2/XIN0/MM0 VREF<0> ENL6<0> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXICDRVP0/XICDRV7/XITIE0/XIN1/MM0 XICDRVP0/XICDRV7/XITIE0/net5 XICDRVP0/XICDRV7/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV7/XITIE0/XIN0/MM0 XICDRVP0/XICDRV7/XITIE0/net6 XICDRVP0/XICDRV7/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXICDRVP0/XICDRV7/XISW0/XIN1/MM0 VREF<2> ENL7<2> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW0/XIN0/MM0 VREF<2> ENL7<2> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW1/XIN1/MM0 VREF<1> ENL7<1> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW1/XIN0/MM0 VREF<1> ENL7<1> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW2/XIN1/MM0 VREF<0> ENL7<0> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXICDRVP0/XICDRV7/XISW2/XIN0/MM0 VREF<0> ENL7<0> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
XICAPM0/XI7<99> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<98> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<97> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<96> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<95> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<94> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<93> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<92> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<91> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<90> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<89> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<88> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<87> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<86> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<85> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<84> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<83> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<82> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<81> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<80> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<79> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<78> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<77> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<76> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<75> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<74> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<73> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<72> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<71> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<70> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<69> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<68> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<67> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<66> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<65> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<64> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<63> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<62> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<61> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<60> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<59> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<58> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<57> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<56> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<55> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<54> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<53> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<52> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<51> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<50> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<49> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<48> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<47> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<46> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<45> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<44> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<43> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<42> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<41> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<40> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<39> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<38> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<37> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<36> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<35> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<34> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<33> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<32> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<31> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<30> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<29> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<28> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<27> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<26> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<25> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<24> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<23> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<22> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<21> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<20> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<19> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<18> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<17> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<16> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<15> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<14> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<13> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<12> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<11> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<10> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<9> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<8> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<7> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<6> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<5> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<4> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<3> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<2> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<1> VOR<7> INM momcap_center_1x 
XICAPM0/XI7<0> VOR<7> INM momcap_center_1x 
XICAPM0/XI6<52> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<51> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<50> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<49> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<48> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<47> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<46> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<45> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<44> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<43> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<42> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<41> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<40> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<39> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<38> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<37> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<36> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<35> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<34> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<33> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<32> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<31> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<30> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<29> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<28> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<27> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<26> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<25> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<24> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<23> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<22> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<21> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<20> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<19> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<18> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<17> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<16> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<15> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<14> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<13> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<12> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<11> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<10> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<9> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<8> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<7> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<6> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<5> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<4> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<3> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<2> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<1> VOR<6> INM momcap_center_1x 
XICAPM0/XI6<0> VOR<6> INM momcap_center_1x 
XICAPM0/XI5<27> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<26> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<25> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<24> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<23> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<22> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<21> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<20> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<19> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<18> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<17> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<16> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<15> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<14> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<13> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<12> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<11> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<10> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<9> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<8> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<7> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<6> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<5> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<4> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<3> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<2> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<1> VOR<5> INM momcap_center_1x 
XICAPM0/XI5<0> VOR<5> INM momcap_center_1x 
XICAPM0/XI4<15> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<14> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<13> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<12> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<11> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<10> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<9> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<8> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<7> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<6> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<5> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<4> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<3> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<2> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<1> VOR<4> INM momcap_center_1x 
XICAPM0/XI4<0> VOR<4> INM momcap_center_1x 
XICAPM0/XI3<7> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<6> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<5> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<4> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<3> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<2> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<1> VOR<3> INM momcap_center_1x 
XICAPM0/XI3<0> VOR<3> INM momcap_center_1x 
XICAPM0/XI2<3> VOR<2> INM momcap_center_1x 
XICAPM0/XI2<2> VOR<2> INM momcap_center_1x 
XICAPM0/XI2<1> VOR<2> INM momcap_center_1x 
XICAPM0/XI2<0> VOR<2> INM momcap_center_1x 
XICAPM0/XI1<1> VOR<1> INM momcap_center_1x 
XICAPM0/XI1<0> VOR<1> INM momcap_center_1x 
XICAPM0/XIC0_0 VREF<1> INM momcap_center_1x 
XICAPM0/XI0 VOR<0> INM momcap_center_1x 
XICAPP0/XI7<99> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<98> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<97> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<96> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<95> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<94> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<93> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<92> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<91> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<90> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<89> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<88> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<87> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<86> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<85> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<84> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<83> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<82> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<81> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<80> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<79> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<78> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<77> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<76> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<75> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<74> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<73> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<72> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<71> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<70> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<69> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<68> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<67> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<66> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<65> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<64> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<63> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<62> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<61> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<60> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<59> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<58> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<57> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<56> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<55> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<54> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<53> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<52> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<51> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<50> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<49> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<48> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<47> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<46> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<45> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<44> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<43> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<42> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<41> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<40> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<39> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<38> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<37> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<36> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<35> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<34> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<33> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<32> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<31> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<30> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<29> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<28> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<27> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<26> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<25> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<24> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<23> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<22> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<21> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<20> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<19> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<18> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<17> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<16> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<15> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<14> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<13> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<12> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<11> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<10> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<9> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<8> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<7> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<6> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<5> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<4> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<3> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<2> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<1> VOL<7> INP momcap_center_1x 
XICAPP0/XI7<0> VOL<7> INP momcap_center_1x 
XICAPP0/XI6<52> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<51> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<50> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<49> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<48> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<47> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<46> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<45> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<44> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<43> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<42> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<41> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<40> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<39> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<38> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<37> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<36> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<35> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<34> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<33> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<32> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<31> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<30> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<29> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<28> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<27> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<26> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<25> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<24> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<23> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<22> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<21> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<20> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<19> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<18> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<17> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<16> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<15> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<14> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<13> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<12> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<11> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<10> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<9> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<8> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<7> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<6> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<5> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<4> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<3> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<2> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<1> VOL<6> INP momcap_center_1x 
XICAPP0/XI6<0> VOL<6> INP momcap_center_1x 
XICAPP0/XI5<27> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<26> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<25> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<24> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<23> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<22> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<21> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<20> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<19> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<18> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<17> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<16> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<15> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<14> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<13> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<12> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<11> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<10> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<9> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<8> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<7> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<6> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<5> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<4> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<3> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<2> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<1> VOL<5> INP momcap_center_1x 
XICAPP0/XI5<0> VOL<5> INP momcap_center_1x 
XICAPP0/XI4<15> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<14> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<13> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<12> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<11> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<10> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<9> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<8> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<7> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<6> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<5> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<4> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<3> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<2> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<1> VOL<4> INP momcap_center_1x 
XICAPP0/XI4<0> VOL<4> INP momcap_center_1x 
XICAPP0/XI3<7> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<6> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<5> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<4> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<3> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<2> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<1> VOL<3> INP momcap_center_1x 
XICAPP0/XI3<0> VOL<3> INP momcap_center_1x 
XICAPP0/XI2<3> VOL<2> INP momcap_center_1x 
XICAPP0/XI2<2> VOL<2> INP momcap_center_1x 
XICAPP0/XI2<1> VOL<2> INP momcap_center_1x 
XICAPP0/XI2<0> VOL<2> INP momcap_center_1x 
XICAPP0/XI1<1> VOL<1> INP momcap_center_1x 
XICAPP0/XI1<0> VOL<1> INP momcap_center_1x 
XICAPP0/XIC0_0 VREF<1> INP momcap_center_1x 
XICAPP0/XI0 VOL<0> INP momcap_center_1x 
.ends

.subckt momcap_center_1x BOTTOM TOP 
.ends

